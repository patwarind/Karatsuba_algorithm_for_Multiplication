`timescale 1ns / 1ps 
//////////////////////////////////////////////////////////////////////////////////  
// Company:    
 // Engineer:   
 //  // Create Date: 25.01.2022 23:34:48 
// Design Name:     
// Module Name: overlap_module 
 // Project Name:    
// Target Devices:  
// Tool Versions:   
// Description: 
//              
// Dependencies:   
 //  
// Revision:       
 // Revision 0.01 - File Created 
// Additional Comments: 
//  
//////////////////////////////////////////////////////////////////////////////////  
    
    
module overlap_module_193bit(     
    B2_in1,                
    B2_in2,             
    B2_in3,   
    B2_out 
    );     


parameter n = 194;
    
input [n-2:0] B2_in1;   
input [n-2:0] B2_in2;    
input [n-2:0] B2_in3;    

output [2*n-2:0] B2_out;  
    


assign B2_out[0] = B2_in1[0];

assign B2_out[1] = B2_in1[1];

assign B2_out[2] = B2_in1[2];

assign B2_out[3] = B2_in1[3];

assign B2_out[4] = B2_in1[4];

assign B2_out[5] = B2_in1[5];

assign B2_out[6] = B2_in1[6];

assign B2_out[7] = B2_in1[7];

assign B2_out[8] = B2_in1[8];

assign B2_out[9] = B2_in1[9];

assign B2_out[10] = B2_in1[10];

assign B2_out[11] = B2_in1[11];

assign B2_out[12] = B2_in1[12];

assign B2_out[13] = B2_in1[13];

assign B2_out[14] = B2_in1[14];

assign B2_out[15] = B2_in1[15];

assign B2_out[16] = B2_in1[16];

assign B2_out[17] = B2_in1[17];

assign B2_out[18] = B2_in1[18];

assign B2_out[19] = B2_in1[19];

assign B2_out[20] = B2_in1[20];

assign B2_out[21] = B2_in1[21];

assign B2_out[22] = B2_in1[22];

assign B2_out[23] = B2_in1[23];

assign B2_out[24] = B2_in1[24];

assign B2_out[25] = B2_in1[25];

assign B2_out[26] = B2_in1[26];

assign B2_out[27] = B2_in1[27];

assign B2_out[28] = B2_in1[28];

assign B2_out[29] = B2_in1[29];

assign B2_out[30] = B2_in1[30];

assign B2_out[31] = B2_in1[31];

assign B2_out[32] = B2_in1[32];

assign B2_out[33] = B2_in1[33];

assign B2_out[34] = B2_in1[34];

assign B2_out[35] = B2_in1[35];

assign B2_out[36] = B2_in1[36];

assign B2_out[37] = B2_in1[37];

assign B2_out[38] = B2_in1[38];

assign B2_out[39] = B2_in1[39];

assign B2_out[40] = B2_in1[40];

assign B2_out[41] = B2_in1[41];

assign B2_out[42] = B2_in1[42];

assign B2_out[43] = B2_in1[43];

assign B2_out[44] = B2_in1[44];

assign B2_out[45] = B2_in1[45];

assign B2_out[46] = B2_in1[46];

assign B2_out[47] = B2_in1[47];

assign B2_out[48] = B2_in1[48];

assign B2_out[49] = B2_in1[49];

assign B2_out[50] = B2_in1[50];

assign B2_out[51] = B2_in1[51];

assign B2_out[52] = B2_in1[52];

assign B2_out[53] = B2_in1[53];

assign B2_out[54] = B2_in1[54];

assign B2_out[55] = B2_in1[55];

assign B2_out[56] = B2_in1[56];

assign B2_out[57] = B2_in1[57];

assign B2_out[58] = B2_in1[58];

assign B2_out[59] = B2_in1[59];

assign B2_out[60] = B2_in1[60];

assign B2_out[61] = B2_in1[61];

assign B2_out[62] = B2_in1[62];

assign B2_out[63] = B2_in1[63];

assign B2_out[64] = B2_in1[64];

assign B2_out[65] = B2_in1[65];

assign B2_out[66] = B2_in1[66];

assign B2_out[67] = B2_in1[67];

assign B2_out[68] = B2_in1[68];

assign B2_out[69] = B2_in1[69];

assign B2_out[70] = B2_in1[70];

assign B2_out[71] = B2_in1[71];

assign B2_out[72] = B2_in1[72];

assign B2_out[73] = B2_in1[73];

assign B2_out[74] = B2_in1[74];

assign B2_out[75] = B2_in1[75];

assign B2_out[76] = B2_in1[76];

assign B2_out[77] = B2_in1[77];

assign B2_out[78] = B2_in1[78];

assign B2_out[79] = B2_in1[79];

assign B2_out[80] = B2_in1[80];

assign B2_out[81] = B2_in1[81];

assign B2_out[82] = B2_in1[82];

assign B2_out[83] = B2_in1[83];

assign B2_out[84] = B2_in1[84];

assign B2_out[85] = B2_in1[85];

assign B2_out[86] = B2_in1[86];

assign B2_out[87] = B2_in1[87];

assign B2_out[88] = B2_in1[88];

assign B2_out[89] = B2_in1[89];

assign B2_out[90] = B2_in1[90];

assign B2_out[91] = B2_in1[91];

assign B2_out[92] = B2_in1[92];

assign B2_out[93] = B2_in1[93];

assign B2_out[94] = B2_in1[94];

assign B2_out[95] = B2_in1[95];

assign B2_out[96] = B2_in1[96];

assign B2_out[97] = B2_in1[97]^ B2_in2[0];

assign B2_out[98] = B2_in1[98]^ B2_in2[1];

assign B2_out[99] = B2_in1[99]^ B2_in2[2];

assign B2_out[100] = B2_in1[100]^ B2_in2[3];

assign B2_out[101] = B2_in1[101]^ B2_in2[4];

assign B2_out[102] = B2_in1[102]^ B2_in2[5];

assign B2_out[103] = B2_in1[103]^ B2_in2[6];

assign B2_out[104] = B2_in1[104]^ B2_in2[7];

assign B2_out[105] = B2_in1[105]^ B2_in2[8];

assign B2_out[106] = B2_in1[106]^ B2_in2[9];

assign B2_out[107] = B2_in1[107]^ B2_in2[10];

assign B2_out[108] = B2_in1[108]^ B2_in2[11];

assign B2_out[109] = B2_in1[109]^ B2_in2[12];

assign B2_out[110] = B2_in1[110]^ B2_in2[13];

assign B2_out[111] = B2_in1[111]^ B2_in2[14];

assign B2_out[112] = B2_in1[112]^ B2_in2[15];

assign B2_out[113] = B2_in1[113]^ B2_in2[16];

assign B2_out[114] = B2_in1[114]^ B2_in2[17];

assign B2_out[115] = B2_in1[115]^ B2_in2[18];

assign B2_out[116] = B2_in1[116]^ B2_in2[19];

assign B2_out[117] = B2_in1[117]^ B2_in2[20];

assign B2_out[118] = B2_in1[118]^ B2_in2[21];

assign B2_out[119] = B2_in1[119]^ B2_in2[22];

assign B2_out[120] = B2_in1[120]^ B2_in2[23];

assign B2_out[121] = B2_in1[121]^ B2_in2[24];

assign B2_out[122] = B2_in1[122]^ B2_in2[25];

assign B2_out[123] = B2_in1[123]^ B2_in2[26];

assign B2_out[124] = B2_in1[124]^ B2_in2[27];

assign B2_out[125] = B2_in1[125]^ B2_in2[28];

assign B2_out[126] = B2_in1[126]^ B2_in2[29];

assign B2_out[127] = B2_in1[127]^ B2_in2[30];

assign B2_out[128] = B2_in1[128]^ B2_in2[31];

assign B2_out[129] = B2_in1[129]^ B2_in2[32];

assign B2_out[130] = B2_in1[130]^ B2_in2[33];

assign B2_out[131] = B2_in1[131]^ B2_in2[34];

assign B2_out[132] = B2_in1[132]^ B2_in2[35];

assign B2_out[133] = B2_in1[133]^ B2_in2[36];

assign B2_out[134] = B2_in1[134]^ B2_in2[37];

assign B2_out[135] = B2_in1[135]^ B2_in2[38];

assign B2_out[136] = B2_in1[136]^ B2_in2[39];

assign B2_out[137] = B2_in1[137]^ B2_in2[40];

assign B2_out[138] = B2_in1[138]^ B2_in2[41];

assign B2_out[139] = B2_in1[139]^ B2_in2[42];

assign B2_out[140] = B2_in1[140]^ B2_in2[43];

assign B2_out[141] = B2_in1[141]^ B2_in2[44];

assign B2_out[142] = B2_in1[142]^ B2_in2[45];

assign B2_out[143] = B2_in1[143]^ B2_in2[46];

assign B2_out[144] = B2_in1[144]^ B2_in2[47];

assign B2_out[145] = B2_in1[145]^ B2_in2[48];

assign B2_out[146] = B2_in1[146]^ B2_in2[49];

assign B2_out[147] = B2_in1[147]^ B2_in2[50];

assign B2_out[148] = B2_in1[148]^ B2_in2[51];

assign B2_out[149] = B2_in1[149]^ B2_in2[52];

assign B2_out[150] = B2_in1[150]^ B2_in2[53];

assign B2_out[151] = B2_in1[151]^ B2_in2[54];

assign B2_out[152] = B2_in1[152]^ B2_in2[55];

assign B2_out[153] = B2_in1[153]^ B2_in2[56];

assign B2_out[154] = B2_in1[154]^ B2_in2[57];

assign B2_out[155] = B2_in1[155]^ B2_in2[58];

assign B2_out[156] = B2_in1[156]^ B2_in2[59];

assign B2_out[157] = B2_in1[157]^ B2_in2[60];

assign B2_out[158] = B2_in1[158]^ B2_in2[61];

assign B2_out[159] = B2_in1[159]^ B2_in2[62];

assign B2_out[160] = B2_in1[160]^ B2_in2[63];

assign B2_out[161] = B2_in1[161]^ B2_in2[64];

assign B2_out[162] = B2_in1[162]^ B2_in2[65];

assign B2_out[163] = B2_in1[163]^ B2_in2[66];

assign B2_out[164] = B2_in1[164]^ B2_in2[67];

assign B2_out[165] = B2_in1[165]^ B2_in2[68];

assign B2_out[166] = B2_in1[166]^ B2_in2[69];

assign B2_out[167] = B2_in1[167]^ B2_in2[70];

assign B2_out[168] = B2_in1[168]^ B2_in2[71];

assign B2_out[169] = B2_in1[169]^ B2_in2[72];

assign B2_out[170] = B2_in1[170]^ B2_in2[73];

assign B2_out[171] = B2_in1[171]^ B2_in2[74];

assign B2_out[172] = B2_in1[172]^ B2_in2[75];

assign B2_out[173] = B2_in1[173]^ B2_in2[76];

assign B2_out[174] = B2_in1[174]^ B2_in2[77];

assign B2_out[175] = B2_in1[175]^ B2_in2[78];

assign B2_out[176] = B2_in1[176]^ B2_in2[79];

assign B2_out[177] = B2_in1[177]^ B2_in2[80];

assign B2_out[178] = B2_in1[178]^ B2_in2[81];

assign B2_out[179] = B2_in1[179]^ B2_in2[82];

assign B2_out[180] = B2_in1[180]^ B2_in2[83];

assign B2_out[181] = B2_in1[181]^ B2_in2[84];

assign B2_out[182] = B2_in1[182]^ B2_in2[85];

assign B2_out[183] = B2_in1[183]^ B2_in2[86];

assign B2_out[184] = B2_in1[184]^ B2_in2[87];

assign B2_out[185] = B2_in1[185]^ B2_in2[88];

assign B2_out[186] = B2_in1[186]^ B2_in2[89];

assign B2_out[187] = B2_in1[187]^ B2_in2[90];

assign B2_out[188] = B2_in1[188]^ B2_in2[91];

assign B2_out[189] = B2_in1[189]^ B2_in2[92];

assign B2_out[190] = B2_in1[190]^ B2_in2[93];

assign B2_out[191] = B2_in1[191]^ B2_in2[94];

assign B2_out[192] = B2_in1[192]^ B2_in2[95];

assign B2_out[193] = B2_in2[96];

assign B2_out[194] = B2_in2[97]^B2_in3[0];

assign B2_out[195] = B2_in2[98]^B2_in3[1];

assign B2_out[196] = B2_in2[99]^B2_in3[2];

assign B2_out[197] = B2_in2[100]^B2_in3[3];

assign B2_out[198] = B2_in2[101]^B2_in3[4];

assign B2_out[199] = B2_in2[102]^B2_in3[5];

assign B2_out[200] = B2_in2[103]^B2_in3[6];

assign B2_out[201] = B2_in2[104]^B2_in3[7];

assign B2_out[202] = B2_in2[105]^B2_in3[8];

assign B2_out[203] = B2_in2[106]^B2_in3[9];

assign B2_out[204] = B2_in2[107]^B2_in3[10];

assign B2_out[205] = B2_in2[108]^B2_in3[11];

assign B2_out[206] = B2_in2[109]^B2_in3[12];

assign B2_out[207] = B2_in2[110]^B2_in3[13];

assign B2_out[208] = B2_in2[111]^B2_in3[14];

assign B2_out[209] = B2_in2[112]^B2_in3[15];

assign B2_out[210] = B2_in2[113]^B2_in3[16];

assign B2_out[211] = B2_in2[114]^B2_in3[17];

assign B2_out[212] = B2_in2[115]^B2_in3[18];

assign B2_out[213] = B2_in2[116]^B2_in3[19];

assign B2_out[214] = B2_in2[117]^B2_in3[20];

assign B2_out[215] = B2_in2[118]^B2_in3[21];

assign B2_out[216] = B2_in2[119]^B2_in3[22];

assign B2_out[217] = B2_in2[120]^B2_in3[23];

assign B2_out[218] = B2_in2[121]^B2_in3[24];

assign B2_out[219] = B2_in2[122]^B2_in3[25];

assign B2_out[220] = B2_in2[123]^B2_in3[26];

assign B2_out[221] = B2_in2[124]^B2_in3[27];

assign B2_out[222] = B2_in2[125]^B2_in3[28];

assign B2_out[223] = B2_in2[126]^B2_in3[29];

assign B2_out[224] = B2_in2[127]^B2_in3[30];

assign B2_out[225] = B2_in2[128]^B2_in3[31];

assign B2_out[226] = B2_in2[129]^B2_in3[32];

assign B2_out[227] = B2_in2[130]^B2_in3[33];

assign B2_out[228] = B2_in2[131]^B2_in3[34];

assign B2_out[229] = B2_in2[132]^B2_in3[35];

assign B2_out[230] = B2_in2[133]^B2_in3[36];

assign B2_out[231] = B2_in2[134]^B2_in3[37];

assign B2_out[232] = B2_in2[135]^B2_in3[38];

assign B2_out[233] = B2_in2[136]^B2_in3[39];

assign B2_out[234] = B2_in2[137]^B2_in3[40];

assign B2_out[235] = B2_in2[138]^B2_in3[41];

assign B2_out[236] = B2_in2[139]^B2_in3[42];

assign B2_out[237] = B2_in2[140]^B2_in3[43];

assign B2_out[238] = B2_in2[141]^B2_in3[44];

assign B2_out[239] = B2_in2[142]^B2_in3[45];

assign B2_out[240] = B2_in2[143]^B2_in3[46];

assign B2_out[241] = B2_in2[144]^B2_in3[47];

assign B2_out[242] = B2_in2[145]^B2_in3[48];

assign B2_out[243] = B2_in2[146]^B2_in3[49];

assign B2_out[244] = B2_in2[147]^B2_in3[50];

assign B2_out[245] = B2_in2[148]^B2_in3[51];

assign B2_out[246] = B2_in2[149]^B2_in3[52];

assign B2_out[247] = B2_in2[150]^B2_in3[53];

assign B2_out[248] = B2_in2[151]^B2_in3[54];

assign B2_out[249] = B2_in2[152]^B2_in3[55];

assign B2_out[250] = B2_in2[153]^B2_in3[56];

assign B2_out[251] = B2_in2[154]^B2_in3[57];

assign B2_out[252] = B2_in2[155]^B2_in3[58];

assign B2_out[253] = B2_in2[156]^B2_in3[59];

assign B2_out[254] = B2_in2[157]^B2_in3[60];

assign B2_out[255] = B2_in2[158]^B2_in3[61];

assign B2_out[256] = B2_in2[159]^B2_in3[62];

assign B2_out[257] = B2_in2[160]^B2_in3[63];

assign B2_out[258] = B2_in2[161]^B2_in3[64];

assign B2_out[259] = B2_in2[162]^B2_in3[65];

assign B2_out[260] = B2_in2[163]^B2_in3[66];

assign B2_out[261] = B2_in2[164]^B2_in3[67];

assign B2_out[262] = B2_in2[165]^B2_in3[68];

assign B2_out[263] = B2_in2[166]^B2_in3[69];

assign B2_out[264] = B2_in2[167]^B2_in3[70];

assign B2_out[265] = B2_in2[168]^B2_in3[71];

assign B2_out[266] = B2_in2[169]^B2_in3[72];

assign B2_out[267] = B2_in2[170]^B2_in3[73];

assign B2_out[268] = B2_in2[171]^B2_in3[74];

assign B2_out[269] = B2_in2[172]^B2_in3[75];

assign B2_out[270] = B2_in2[173]^B2_in3[76];

assign B2_out[271] = B2_in2[174]^B2_in3[77];

assign B2_out[272] = B2_in2[175]^B2_in3[78];

assign B2_out[273] = B2_in2[176]^B2_in3[79];

assign B2_out[274] = B2_in2[177]^B2_in3[80];

assign B2_out[275] = B2_in2[178]^B2_in3[81];

assign B2_out[276] = B2_in2[179]^B2_in3[82];

assign B2_out[277] = B2_in2[180]^B2_in3[83];

assign B2_out[278] = B2_in2[181]^B2_in3[84];

assign B2_out[279] = B2_in2[182]^B2_in3[85];

assign B2_out[280] = B2_in2[183]^B2_in3[86];

assign B2_out[281] = B2_in2[184]^B2_in3[87];

assign B2_out[282] = B2_in2[185]^B2_in3[88];

assign B2_out[283] = B2_in2[186]^B2_in3[89];

assign B2_out[284] = B2_in2[187]^B2_in3[90];

assign B2_out[285] = B2_in2[188]^B2_in3[91];

assign B2_out[286] = B2_in2[189]^B2_in3[92];

assign B2_out[287] = B2_in2[190]^B2_in3[93];

assign B2_out[288] = B2_in2[191]^B2_in3[94];

assign B2_out[289] = B2_in2[192]^B2_in3[95];

assign B2_out[290] = B2_in3[96];

assign B2_out[291] = B2_in3[97];

assign B2_out[292] = B2_in3[98];

assign B2_out[293] = B2_in3[99];

assign B2_out[294] = B2_in3[100];

assign B2_out[295] = B2_in3[101];

assign B2_out[296] = B2_in3[102];

assign B2_out[297] = B2_in3[103];

assign B2_out[298] = B2_in3[104];

assign B2_out[299] = B2_in3[105];

assign B2_out[300] = B2_in3[106];

assign B2_out[301] = B2_in3[107];

assign B2_out[302] = B2_in3[108];

assign B2_out[303] = B2_in3[109];

assign B2_out[304] = B2_in3[110];

assign B2_out[305] = B2_in3[111];

assign B2_out[306] = B2_in3[112];

assign B2_out[307] = B2_in3[113];

assign B2_out[308] = B2_in3[114];

assign B2_out[309] = B2_in3[115];

assign B2_out[310] = B2_in3[116];

assign B2_out[311] = B2_in3[117];

assign B2_out[312] = B2_in3[118];

assign B2_out[313] = B2_in3[119];

assign B2_out[314] = B2_in3[120];

assign B2_out[315] = B2_in3[121];

assign B2_out[316] = B2_in3[122];

assign B2_out[317] = B2_in3[123];

assign B2_out[318] = B2_in3[124];

assign B2_out[319] = B2_in3[125];

assign B2_out[320] = B2_in3[126];

assign B2_out[321] = B2_in3[127];

assign B2_out[322] = B2_in3[128];

assign B2_out[323] = B2_in3[129];

assign B2_out[324] = B2_in3[130];

assign B2_out[325] = B2_in3[131];

assign B2_out[326] = B2_in3[132];

assign B2_out[327] = B2_in3[133];

assign B2_out[328] = B2_in3[134];

assign B2_out[329] = B2_in3[135];

assign B2_out[330] = B2_in3[136];

assign B2_out[331] = B2_in3[137];

assign B2_out[332] = B2_in3[138];

assign B2_out[333] = B2_in3[139];

assign B2_out[334] = B2_in3[140];

assign B2_out[335] = B2_in3[141];

assign B2_out[336] = B2_in3[142];

assign B2_out[337] = B2_in3[143];

assign B2_out[338] = B2_in3[144];

assign B2_out[339] = B2_in3[145];

assign B2_out[340] = B2_in3[146];

assign B2_out[341] = B2_in3[147];

assign B2_out[342] = B2_in3[148];

assign B2_out[343] = B2_in3[149];

assign B2_out[344] = B2_in3[150];

assign B2_out[345] = B2_in3[151];

assign B2_out[346] = B2_in3[152];

assign B2_out[347] = B2_in3[153];

assign B2_out[348] = B2_in3[154];

assign B2_out[349] = B2_in3[155];

assign B2_out[350] = B2_in3[156];

assign B2_out[351] = B2_in3[157];

assign B2_out[352] = B2_in3[158];

assign B2_out[353] = B2_in3[159];

assign B2_out[354] = B2_in3[160];

assign B2_out[355] = B2_in3[161];

assign B2_out[356] = B2_in3[162];

assign B2_out[357] = B2_in3[163];

assign B2_out[358] = B2_in3[164];

assign B2_out[359] = B2_in3[165];

assign B2_out[360] = B2_in3[166];

assign B2_out[361] = B2_in3[167];

assign B2_out[362] = B2_in3[168];

assign B2_out[363] = B2_in3[169];

assign B2_out[364] = B2_in3[170];

assign B2_out[365] = B2_in3[171];

assign B2_out[366] = B2_in3[172];

assign B2_out[367] = B2_in3[173];

assign B2_out[368] = B2_in3[174];

assign B2_out[369] = B2_in3[175];

assign B2_out[370] = B2_in3[176];

assign B2_out[371] = B2_in3[177];

assign B2_out[372] = B2_in3[178];

assign B2_out[373] = B2_in3[179];

assign B2_out[374] = B2_in3[180];

assign B2_out[375] = B2_in3[181];

assign B2_out[376] = B2_in3[182];

assign B2_out[377] = B2_in3[183];

assign B2_out[378] = B2_in3[184];

assign B2_out[379] = B2_in3[185];

assign B2_out[380] = B2_in3[186];

assign B2_out[381] = B2_in3[187];

assign B2_out[382] = B2_in3[188];

assign B2_out[383] = B2_in3[189];

assign B2_out[384] = B2_in3[190];

assign B2_out[385] = B2_in3[191];

assign B2_out[386] = B2_in3[192];

endmodule